module INST_MEM(
    clk,
    reset,
    read_address,
    instruction_out
);

input clk, reset;
input [31:0] read_address;
output [31:0] instruction_out;
reg [31:0] I_Mem[63:0];
//integer k;
assign instruction_out = I_Mem[read_address];
/*initial begin
    I_Mem[0]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[1]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[2]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[3]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[4]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[5]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[6]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[7]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[8]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[9]  <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[10] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[11] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[12] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[13] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[14] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[15] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[16] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[17] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[18] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[19] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[20] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[21] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[22] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[23] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[24] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[25] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[26] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[27] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[28] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[29] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[30] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[31] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[32] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[33] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[34] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[35] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[36] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[37] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[38] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[39] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[40] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[41] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[42] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[43] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[44] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[45] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[46] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[47] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[48] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[49] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[50] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[51] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[52] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[53] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[54] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[55] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[56] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[57] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[58] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[59] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[60] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[61] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[62] <= 32'b0000000_00000_00000_000_00000_0000000;
    I_Mem[63] <= 32'b0000000_00000_00000_000_00000_0000000;
end
*/

always @(posedge clk or posedge reset)
begin

if(reset)
    begin   
        /*for(k=0;k<64;k=k+1) begin
        I_Mem[k] <= 32'b00;
        end */
        
        //I_Mem[0] <= 32'b0000000_00000_00000_000_00000_0000000; // no operation
         I_Mem[0]  <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[1]  <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[2]  <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[3]  <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[4]  <= 32'b0000000_11001_10000_000_01101_0110011; // add x13, x16, x25
           I_Mem[5]  <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[6]  <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[7]  <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[8]  <= 32'b0100000_00011_01000_000_00101_0110011; // sub x5, x8, x3
           I_Mem[9]  <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[10] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[11] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[12] <= 32'b0000000_00011_00010_111_00001_0110011;// and x1, x2, x3
           I_Mem[13] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[14] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[15] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[16] <= 32'b0000000_00101_00011_110_00100_0110011; // or x4, x3, x5
           I_Mem[17] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[18] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[19] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[20] <= 32'b000000000011_10101_000_10110_0010011; // addi x22, x21, 3
           I_Mem[21] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[22] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[23] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[24] <= 32'b000000000001_01000_110_01001_0010011; // ori x9, x8, 1
           I_Mem[25] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[26] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[27] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[28] <= 32'b000000001111_00101_010_01000_0000011; // lw x8, 15(x5)
           I_Mem[29] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[30] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[31] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[32] <= 32'b000000000011_00011_010_01001_0000011; // lw x9, 3(x3)
           I_Mem[33] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[34] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[35] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[36] <= 32'b0000000_01111_00101_010_01100_0100011;// sw x15, 12(x5)
           I_Mem[37] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[38] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[39] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[40] <= 32'b0000000_01110_00110_010_01010_0100011;// sw x14, 10(x6)
           I_Mem[41] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[42] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[43] <= 32'b0000000_00000_00000_000_00000_0000000;
           //I_Mem[44] <= 32'h00948663; // beq x9, x9, 12
           I_Mem[44] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[45] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[46] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[47] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[48] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[49] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[50] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[51] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[52] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[53] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[54] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[55] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[56] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[57] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[58] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[59] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[60] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[61] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[62] <= 32'b0000000_00000_00000_000_00000_0000000;
           I_Mem[63] <= 32'b0000000_00000_00000_000_00000_0000000;
                
    end
//else

   //I_Mem[0] = 32'b0000000_00000_00000_000_00000_0000000; // no operation
   
 /*
    // R-Type
        I_Mem[4] = 32'b0000000_11001_10000_000_01101_0110011; // add x13, x16, x25
        I_Mem[8] = 32'b0100000_00011_01000_000_00101_0110011; // sub x5, x8, x3
        I_Mem[12] = 32'b0000000_00011_00010_111_00001_0110011;// and x1, x2, x3
        I_Mem[16] = 32'b0000000_00101_00011_110_00100_0110011; // or x4, x3, x5

    // I-Type
        I_Mem[20] = 32'b000000000011_10101_000_10110_0010011; // addi x22, x21, 3
        I_Mem[24] = 32'b000000000001_01000_110_01001_0010011; // ori x9, x8, 1

    // L-Type
        I_Mem[28] = 32'b000000001111_00101_010_01000_0000011; // lw x8, 15(x5)
        I_Mem[32] = 32'b000000000011_00011_010_01001_0000011; // lw x9, 3(x3)
    
    // S-Type
        I_Mem[36] = 32'b0000000_01111_00101_010_01100_0100011;// sw x15, 12(x5)
        I_Mem[40] = 32'b0000000_01110_00110_010_01010_0100011;// sw x14, 10(x6)
    
    // SB-Type
        I_Mem[44] = 32'h00948663; // beq x9, x9, 12 */

end
endmodule
